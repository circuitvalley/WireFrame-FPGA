library verilog;
use verilog.vl_types.all;
entity counter_testbench is
end counter_testbench;
